module ast

pub interface Node {
	display()
}
