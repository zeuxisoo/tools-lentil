module expressions

pub struct IdentifierExpression {
	value string
}

pub fn (s IdentifierExpression) display() {
	println('TODO: identifier')
}
