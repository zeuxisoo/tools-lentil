module expressions

pub struct AccountExpression {
mut:
	value string
	kind  string
}

pub fn (a AccountExpression) display() {
	println('TODO: account')
}
