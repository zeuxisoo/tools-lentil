module expressions

import ast { Expression }

pub struct DateRecordsExpression {
pub:
	values []Expression
}

pub fn (dr DateRecordsExpression) display() {
	println('TODO: date records')
}
