module ast

pub interface Expression {
	Node
}
