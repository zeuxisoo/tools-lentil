module ast

pub struct Program {
pub mut:
	statements []Statement
}

fn (p Program) display() {
	println('TODO: Program')
}
