module ast

pub interface Node {
	str() string
}
