module statements

import ast { Statement }

pub struct DateStatement {
	block Statement
}

pub fn (ds DateStatement) display() {
	println('TODO: date statement')
}
