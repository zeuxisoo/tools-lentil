module ast

pub interface Statement {
	Node
}
