module expressions

import ast { Expression }

pub struct AmountsExpression {
	values []Expression
}

pub fn (a AmountsExpression) display() {
	println('TODO: amounts')
}
