module expressions

import ast { Expression }

pub struct DateRecordsExpression {
pub:
	values []Expression
}

pub fn (dr DateRecordsExpression) str() string {
	return 'TODO: date records'
}
