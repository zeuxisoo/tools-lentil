module expressions

pub type Expression = AccountExpression
	| AmountExpression
	| AmountsExpression
	| ArrayExpression
	| AssignExpression
	| AtomExpression
	| DateRecordReceiptExpression
	| DateRecordExpression
	| DateRecordsExpression
	| IdentifierExpression
	| NumberKindExpression
	| NumberExpression
	| StringExpression
