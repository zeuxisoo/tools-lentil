module ast

pub interface Statement {
	str() string
}
