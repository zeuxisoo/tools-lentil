module statements

import ast { Expression }

pub struct DateBlockStatement {
	value []Expression
}

pub fn (db DateBlockStatement) display() {
	println('TODO: date block')
}
