module expressions

import ast { Expression }

pub struct AmountsExpression {
pub:
	values []Expression
}

pub fn (a AmountsExpression) str() string {
	return 'TODO: amounts'
}
