module expressions

import ast { Expression }

pub struct NumberKindExpression {
	value string
}

pub fn (n NumberKindExpression) display() {
	println('TODO: number kind')
}
