module expressions

pub struct NumberKindExpression {
pub:
	value string
}

pub fn (n NumberKindExpression) display() {
	println('TODO: number kind')
}
