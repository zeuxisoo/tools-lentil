module statements

pub struct ConfigStatement {
pub:
	block Statement
}

pub fn (c ConfigStatement) str() string {
	return 'TODO: config'
}
