module expressions

pub struct NumberKindExpression {
	value string
}

pub fn (n NumberKindExpression) display() {
	println('TODO: number kind')
}
