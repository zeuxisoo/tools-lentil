module ast

pub interface Statement {
	display()
}
