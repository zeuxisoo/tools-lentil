module expressions

pub struct AtomExpression {
	value string
}

pub fn (t AtomExpression) display() {
	println('TODO: atom')
}
