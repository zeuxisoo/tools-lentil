module parser

import ast { Expression }
import ast.expressions { DateRecordExpression }

fn parse_date_record_expression(mut parser Parser) !Expression {
	mut expressions := [
		parse_date_record_receipt_expression(mut parser)!
	]

	for parser.current_token.kind in [.bit_wise_and] {
		if parser.current_token.kind == .bit_wise_and {
			parser.read_token()
		}

		expressions << parse_date_record_receipt_expression(mut parser)!
	}

	expression := DateRecordExpression{
		values: expressions
	}

	return expression
}
