module ast

pub interface Expression {
	str() string
}
