module expressions

pub struct AtomExpression {
pub:
	value string
}

pub fn (t AtomExpression) display() {
	println('TODO: atom')
}
