module expressions

pub struct IdentifierExpression {
pub:
	value string
}

pub fn (s IdentifierExpression) str() string {
	return s.value
}
