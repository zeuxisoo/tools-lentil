module expressions

pub struct IdentifierExpression {
pub:
	value string
}

pub fn (s IdentifierExpression) ast() string {
	return s.value
}
