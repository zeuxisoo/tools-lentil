module expressions

import ast { Expression }

pub struct DateRecordExpression {
	values []Expression
}

pub fn (dr DateRecordExpression) display() {
	println('TODO: date record')
}
