module statements

import ast { Statement }

pub struct ConfigStatement {
pub:
	block Statement
}

pub fn (c ConfigStatement) display() {
	println('TODO: config')
}
