module ast

pub interface Expression {
	display()
}
