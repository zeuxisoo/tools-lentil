module expressions

pub struct StringExpression {
pub mut:
	value string
}

pub fn (s StringExpression) display() {
	println('TODO: string')
}
