module expressions

pub struct AccountExpression {
pub mut:
	value string
mut:
	kind  string
}

pub fn (a AccountExpression) display() {
	println('TODO: account')
}
