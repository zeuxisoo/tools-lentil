module expressions

pub struct StringExpression {
mut:
	value string
}

pub fn (s StringExpression) display() {
	println('TODO: string')
}
