module expressions

pub struct IdentifierExpression {
pub:
	value string
}

pub fn (s IdentifierExpression) display() {
	println('TODO: identifier')
}
